// Mk8_Observer_CPU.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module Mk8_Observer_CPU (
		input  wire        altpll_sys_areset_conduit_export,                   //               altpll_sys_areset_conduit.export
		output wire        altpll_sys_locked_conduit_export,                   //               altpll_sys_locked_conduit.export
		input  wire        clk_clk,                                            //                                     clk.clk
		output wire        clk_100m_clk,                                       //                                clk_100m.clk
		output wire        clk_200m_clk,                                       //                                clk_200m.clk
		output wire        cpu_clk_clk,                                        //                                 cpu_clk.clk
		input  wire        external_bus_bridge_external_interface_acknowledge, //  external_bus_bridge_external_interface.acknowledge
		input  wire        external_bus_bridge_external_interface_irq,         //                                        .irq
		output wire [7:0]  external_bus_bridge_external_interface_address,     //                                        .address
		output wire        external_bus_bridge_external_interface_bus_enable,  //                                        .bus_enable
		output wire        external_bus_bridge_external_interface_byte_enable, //                                        .byte_enable
		output wire        external_bus_bridge_external_interface_rw,          //                                        .rw
		output wire [7:0]  external_bus_bridge_external_interface_write_data,  //                                        .write_data
		input  wire [7:0]  external_bus_bridge_external_interface_read_data,   //                                        .read_data
		input  wire        parameter_clk_1_clk,                                //                         parameter_clk_1.clk
		input  wire        parameter_sys_parameter_loop_gpio_in_port,          //       parameter_sys_parameter_loop_gpio.in_port
		output wire        parameter_sys_parameter_loop_gpio_out_port,         //                                        .out_port
		input  wire [10:0] parameter_sys_parameter_rx_ram_s2_address,          //       parameter_sys_parameter_rx_ram_s2.address
		input  wire        parameter_sys_parameter_rx_ram_s2_chipselect,       //                                        .chipselect
		input  wire        parameter_sys_parameter_rx_ram_s2_clken,            //                                        .clken
		input  wire        parameter_sys_parameter_rx_ram_s2_write,            //                                        .write
		output wire [31:0] parameter_sys_parameter_rx_ram_s2_readdata,         //                                        .readdata
		input  wire [31:0] parameter_sys_parameter_rx_ram_s2_writedata,        //                                        .writedata
		input  wire [3:0]  parameter_sys_parameter_rx_ram_s2_byteenable,       //                                        .byteenable
		input  wire [10:0] parameter_sys_parameter_tx_ram_s2_address,          //       parameter_sys_parameter_tx_ram_s2.address
		input  wire        parameter_sys_parameter_tx_ram_s2_chipselect,       //                                        .chipselect
		input  wire        parameter_sys_parameter_tx_ram_s2_clken,            //                                        .clken
		input  wire        parameter_sys_parameter_tx_ram_s2_write,            //                                        .write
		output wire [31:0] parameter_sys_parameter_tx_ram_s2_readdata,         //                                        .readdata
		input  wire [31:0] parameter_sys_parameter_tx_ram_s2_writedata,        //                                        .writedata
		input  wire [3:0]  parameter_sys_parameter_tx_ram_s2_byteenable,       //                                        .byteenable
		output wire        parameter_sys_reset_out_export,                     //                 parameter_sys_reset_out.export
		output wire [7:0]  pheriphals_led_gpio_external_connection_export,     // pheriphals_led_gpio_external_connection.export
		output wire [7:0]  pheriphals_tp_gpio_external_connection_export,      //  pheriphals_tp_gpio_external_connection.export
		input  wire        reset_reset_n,                                      //                                   reset.reset_n
		input  wire        reset_parameter_reset_n                             //                         reset_parameter.reset_n
	);

	wire          vic_0_interrupt_controller_out_valid;                           // vic_0:interrupt_controller_out_valid -> nios2_gen2:eic_port_valid
	wire   [44:0] vic_0_interrupt_controller_out_data;                            // vic_0:interrupt_controller_out_data -> nios2_gen2:eic_port_data
	wire   [31:0] nios2_gen2_data_master_readdata;                                // mm_interconnect_0:nios2_gen2_data_master_readdata -> nios2_gen2:d_readdata
	wire          nios2_gen2_data_master_waitrequest;                             // mm_interconnect_0:nios2_gen2_data_master_waitrequest -> nios2_gen2:d_waitrequest
	wire          nios2_gen2_data_master_debugaccess;                             // nios2_gen2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_data_master_debugaccess
	wire   [18:0] nios2_gen2_data_master_address;                                 // nios2_gen2:d_address -> mm_interconnect_0:nios2_gen2_data_master_address
	wire    [3:0] nios2_gen2_data_master_byteenable;                              // nios2_gen2:d_byteenable -> mm_interconnect_0:nios2_gen2_data_master_byteenable
	wire          nios2_gen2_data_master_read;                                    // nios2_gen2:d_read -> mm_interconnect_0:nios2_gen2_data_master_read
	wire          nios2_gen2_data_master_readdatavalid;                           // mm_interconnect_0:nios2_gen2_data_master_readdatavalid -> nios2_gen2:d_readdatavalid
	wire          nios2_gen2_data_master_write;                                   // nios2_gen2:d_write -> mm_interconnect_0:nios2_gen2_data_master_write
	wire   [31:0] nios2_gen2_data_master_writedata;                               // nios2_gen2:d_writedata -> mm_interconnect_0:nios2_gen2_data_master_writedata
	wire   [31:0] msgdma_0_mm_read_readdata;                                      // mm_interconnect_0:msgdma_0_mm_read_readdata -> msgdma_0:mm_read_readdata
	wire          msgdma_0_mm_read_waitrequest;                                   // mm_interconnect_0:msgdma_0_mm_read_waitrequest -> msgdma_0:mm_read_waitrequest
	wire   [18:0] msgdma_0_mm_read_address;                                       // msgdma_0:mm_read_address -> mm_interconnect_0:msgdma_0_mm_read_address
	wire          msgdma_0_mm_read_read;                                          // msgdma_0:mm_read_read -> mm_interconnect_0:msgdma_0_mm_read_read
	wire    [3:0] msgdma_0_mm_read_byteenable;                                    // msgdma_0:mm_read_byteenable -> mm_interconnect_0:msgdma_0_mm_read_byteenable
	wire          msgdma_0_mm_read_readdatavalid;                                 // mm_interconnect_0:msgdma_0_mm_read_readdatavalid -> msgdma_0:mm_read_readdatavalid
	wire          msgdma_0_mm_write_waitrequest;                                  // mm_interconnect_0:msgdma_0_mm_write_waitrequest -> msgdma_0:mm_write_waitrequest
	wire   [18:0] msgdma_0_mm_write_address;                                      // msgdma_0:mm_write_address -> mm_interconnect_0:msgdma_0_mm_write_address
	wire    [3:0] msgdma_0_mm_write_byteenable;                                   // msgdma_0:mm_write_byteenable -> mm_interconnect_0:msgdma_0_mm_write_byteenable
	wire          msgdma_0_mm_write_write;                                        // msgdma_0:mm_write_write -> mm_interconnect_0:msgdma_0_mm_write_write
	wire   [31:0] msgdma_0_mm_write_writedata;                                    // msgdma_0:mm_write_writedata -> mm_interconnect_0:msgdma_0_mm_write_writedata
	wire   [31:0] nios2_gen2_instruction_master_readdata;                         // mm_interconnect_0:nios2_gen2_instruction_master_readdata -> nios2_gen2:i_readdata
	wire          nios2_gen2_instruction_master_waitrequest;                      // mm_interconnect_0:nios2_gen2_instruction_master_waitrequest -> nios2_gen2:i_waitrequest
	wire   [18:0] nios2_gen2_instruction_master_address;                          // nios2_gen2:i_address -> mm_interconnect_0:nios2_gen2_instruction_master_address
	wire          nios2_gen2_instruction_master_read;                             // nios2_gen2:i_read -> mm_interconnect_0:nios2_gen2_instruction_master_read
	wire          nios2_gen2_instruction_master_readdatavalid;                    // mm_interconnect_0:nios2_gen2_instruction_master_readdatavalid -> nios2_gen2:i_readdatavalid
	wire          mm_interconnect_0_external_bus_bridge_avalon_slave_chipselect;  // mm_interconnect_0:external_bus_bridge_avalon_slave_chipselect -> external_bus_bridge:avalon_chipselect
	wire    [7:0] mm_interconnect_0_external_bus_bridge_avalon_slave_readdata;    // external_bus_bridge:avalon_readdata -> mm_interconnect_0:external_bus_bridge_avalon_slave_readdata
	wire          mm_interconnect_0_external_bus_bridge_avalon_slave_waitrequest; // external_bus_bridge:avalon_waitrequest -> mm_interconnect_0:external_bus_bridge_avalon_slave_waitrequest
	wire    [7:0] mm_interconnect_0_external_bus_bridge_avalon_slave_address;     // mm_interconnect_0:external_bus_bridge_avalon_slave_address -> external_bus_bridge:avalon_address
	wire          mm_interconnect_0_external_bus_bridge_avalon_slave_read;        // mm_interconnect_0:external_bus_bridge_avalon_slave_read -> external_bus_bridge:avalon_read
	wire    [0:0] mm_interconnect_0_external_bus_bridge_avalon_slave_byteenable;  // mm_interconnect_0:external_bus_bridge_avalon_slave_byteenable -> external_bus_bridge:avalon_byteenable
	wire          mm_interconnect_0_external_bus_bridge_avalon_slave_write;       // mm_interconnect_0:external_bus_bridge_avalon_slave_write -> external_bus_bridge:avalon_write
	wire    [7:0] mm_interconnect_0_external_bus_bridge_avalon_slave_writedata;   // mm_interconnect_0:external_bus_bridge_avalon_slave_writedata -> external_bus_bridge:avalon_writedata
	wire   [31:0] mm_interconnect_0_msgdma_0_csr_readdata;                        // msgdma_0:csr_readdata -> mm_interconnect_0:msgdma_0_csr_readdata
	wire    [2:0] mm_interconnect_0_msgdma_0_csr_address;                         // mm_interconnect_0:msgdma_0_csr_address -> msgdma_0:csr_address
	wire          mm_interconnect_0_msgdma_0_csr_read;                            // mm_interconnect_0:msgdma_0_csr_read -> msgdma_0:csr_read
	wire    [3:0] mm_interconnect_0_msgdma_0_csr_byteenable;                      // mm_interconnect_0:msgdma_0_csr_byteenable -> msgdma_0:csr_byteenable
	wire          mm_interconnect_0_msgdma_0_csr_write;                           // mm_interconnect_0:msgdma_0_csr_write -> msgdma_0:csr_write
	wire   [31:0] mm_interconnect_0_msgdma_0_csr_writedata;                       // mm_interconnect_0:msgdma_0_csr_writedata -> msgdma_0:csr_writedata
	wire   [31:0] mm_interconnect_0_vic_0_csr_access_readdata;                    // vic_0:csr_access_readdata -> mm_interconnect_0:vic_0_csr_access_readdata
	wire    [7:0] mm_interconnect_0_vic_0_csr_access_address;                     // mm_interconnect_0:vic_0_csr_access_address -> vic_0:csr_access_address
	wire          mm_interconnect_0_vic_0_csr_access_read;                        // mm_interconnect_0:vic_0_csr_access_read -> vic_0:csr_access_read
	wire          mm_interconnect_0_vic_0_csr_access_write;                       // mm_interconnect_0:vic_0_csr_access_write -> vic_0:csr_access_write
	wire   [31:0] mm_interconnect_0_vic_0_csr_access_writedata;                   // mm_interconnect_0:vic_0_csr_access_writedata -> vic_0:csr_access_writedata
	wire   [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata;          // nios2_gen2:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_debug_mem_slave_readdata
	wire          mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest;       // nios2_gen2:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_debug_mem_slave_waitrequest
	wire          mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess;       // mm_interconnect_0:nios2_gen2_debug_mem_slave_debugaccess -> nios2_gen2:debug_mem_slave_debugaccess
	wire    [8:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_address;           // mm_interconnect_0:nios2_gen2_debug_mem_slave_address -> nios2_gen2:debug_mem_slave_address
	wire          mm_interconnect_0_nios2_gen2_debug_mem_slave_read;              // mm_interconnect_0:nios2_gen2_debug_mem_slave_read -> nios2_gen2:debug_mem_slave_read
	wire    [3:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable;        // mm_interconnect_0:nios2_gen2_debug_mem_slave_byteenable -> nios2_gen2:debug_mem_slave_byteenable
	wire          mm_interconnect_0_nios2_gen2_debug_mem_slave_write;             // mm_interconnect_0:nios2_gen2_debug_mem_slave_write -> nios2_gen2:debug_mem_slave_write
	wire   [31:0] mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata;         // mm_interconnect_0:nios2_gen2_debug_mem_slave_writedata -> nios2_gen2:debug_mem_slave_writedata
	wire          mm_interconnect_0_msgdma_0_descriptor_slave_waitrequest;        // msgdma_0:descriptor_slave_waitrequest -> mm_interconnect_0:msgdma_0_descriptor_slave_waitrequest
	wire   [31:0] mm_interconnect_0_msgdma_0_descriptor_slave_byteenable;         // mm_interconnect_0:msgdma_0_descriptor_slave_byteenable -> msgdma_0:descriptor_slave_byteenable
	wire          mm_interconnect_0_msgdma_0_descriptor_slave_write;              // mm_interconnect_0:msgdma_0_descriptor_slave_write -> msgdma_0:descriptor_slave_write
	wire  [255:0] mm_interconnect_0_msgdma_0_descriptor_slave_writedata;          // mm_interconnect_0:msgdma_0_descriptor_slave_writedata -> msgdma_0:descriptor_slave_writedata
	wire   [31:0] mm_interconnect_0_pheriphals_mapped_slave_readdata;             // Pheriphals:mapped_slave_readdata -> mm_interconnect_0:Pheriphals_mapped_slave_readdata
	wire          mm_interconnect_0_pheriphals_mapped_slave_waitrequest;          // Pheriphals:mapped_slave_waitrequest -> mm_interconnect_0:Pheriphals_mapped_slave_waitrequest
	wire          mm_interconnect_0_pheriphals_mapped_slave_debugaccess;          // mm_interconnect_0:Pheriphals_mapped_slave_debugaccess -> Pheriphals:mapped_slave_debugaccess
	wire    [9:0] mm_interconnect_0_pheriphals_mapped_slave_address;              // mm_interconnect_0:Pheriphals_mapped_slave_address -> Pheriphals:mapped_slave_address
	wire          mm_interconnect_0_pheriphals_mapped_slave_read;                 // mm_interconnect_0:Pheriphals_mapped_slave_read -> Pheriphals:mapped_slave_read
	wire    [3:0] mm_interconnect_0_pheriphals_mapped_slave_byteenable;           // mm_interconnect_0:Pheriphals_mapped_slave_byteenable -> Pheriphals:mapped_slave_byteenable
	wire          mm_interconnect_0_pheriphals_mapped_slave_readdatavalid;        // Pheriphals:mapped_slave_readdatavalid -> mm_interconnect_0:Pheriphals_mapped_slave_readdatavalid
	wire          mm_interconnect_0_pheriphals_mapped_slave_write;                // mm_interconnect_0:Pheriphals_mapped_slave_write -> Pheriphals:mapped_slave_write
	wire   [31:0] mm_interconnect_0_pheriphals_mapped_slave_writedata;            // mm_interconnect_0:Pheriphals_mapped_slave_writedata -> Pheriphals:mapped_slave_writedata
	wire    [0:0] mm_interconnect_0_pheriphals_mapped_slave_burstcount;           // mm_interconnect_0:Pheriphals_mapped_slave_burstcount -> Pheriphals:mapped_slave_burstcount
	wire   [31:0] mm_interconnect_0_timersys_0_mapped_slave_readdata;             // TimerSYS_0:mapped_slave_readdata -> mm_interconnect_0:TimerSYS_0_mapped_slave_readdata
	wire          mm_interconnect_0_timersys_0_mapped_slave_waitrequest;          // TimerSYS_0:mapped_slave_waitrequest -> mm_interconnect_0:TimerSYS_0_mapped_slave_waitrequest
	wire          mm_interconnect_0_timersys_0_mapped_slave_debugaccess;          // mm_interconnect_0:TimerSYS_0_mapped_slave_debugaccess -> TimerSYS_0:mapped_slave_debugaccess
	wire    [9:0] mm_interconnect_0_timersys_0_mapped_slave_address;              // mm_interconnect_0:TimerSYS_0_mapped_slave_address -> TimerSYS_0:mapped_slave_address
	wire          mm_interconnect_0_timersys_0_mapped_slave_read;                 // mm_interconnect_0:TimerSYS_0_mapped_slave_read -> TimerSYS_0:mapped_slave_read
	wire    [3:0] mm_interconnect_0_timersys_0_mapped_slave_byteenable;           // mm_interconnect_0:TimerSYS_0_mapped_slave_byteenable -> TimerSYS_0:mapped_slave_byteenable
	wire          mm_interconnect_0_timersys_0_mapped_slave_readdatavalid;        // TimerSYS_0:mapped_slave_readdatavalid -> mm_interconnect_0:TimerSYS_0_mapped_slave_readdatavalid
	wire          mm_interconnect_0_timersys_0_mapped_slave_write;                // mm_interconnect_0:TimerSYS_0_mapped_slave_write -> TimerSYS_0:mapped_slave_write
	wire   [31:0] mm_interconnect_0_timersys_0_mapped_slave_writedata;            // mm_interconnect_0:TimerSYS_0_mapped_slave_writedata -> TimerSYS_0:mapped_slave_writedata
	wire    [0:0] mm_interconnect_0_timersys_0_mapped_slave_burstcount;           // mm_interconnect_0:TimerSYS_0_mapped_slave_burstcount -> TimerSYS_0:mapped_slave_burstcount
	wire   [31:0] mm_interconnect_0_parameter_sys_mapped_slave_readdata;          // Parameter_SYS:mapped_slave_readdata -> mm_interconnect_0:Parameter_SYS_mapped_slave_readdata
	wire          mm_interconnect_0_parameter_sys_mapped_slave_waitrequest;       // Parameter_SYS:mapped_slave_waitrequest -> mm_interconnect_0:Parameter_SYS_mapped_slave_waitrequest
	wire          mm_interconnect_0_parameter_sys_mapped_slave_debugaccess;       // mm_interconnect_0:Parameter_SYS_mapped_slave_debugaccess -> Parameter_SYS:mapped_slave_debugaccess
	wire   [14:0] mm_interconnect_0_parameter_sys_mapped_slave_address;           // mm_interconnect_0:Parameter_SYS_mapped_slave_address -> Parameter_SYS:mapped_slave_address
	wire          mm_interconnect_0_parameter_sys_mapped_slave_read;              // mm_interconnect_0:Parameter_SYS_mapped_slave_read -> Parameter_SYS:mapped_slave_read
	wire    [3:0] mm_interconnect_0_parameter_sys_mapped_slave_byteenable;        // mm_interconnect_0:Parameter_SYS_mapped_slave_byteenable -> Parameter_SYS:mapped_slave_byteenable
	wire          mm_interconnect_0_parameter_sys_mapped_slave_readdatavalid;     // Parameter_SYS:mapped_slave_readdatavalid -> mm_interconnect_0:Parameter_SYS_mapped_slave_readdatavalid
	wire          mm_interconnect_0_parameter_sys_mapped_slave_write;             // mm_interconnect_0:Parameter_SYS_mapped_slave_write -> Parameter_SYS:mapped_slave_write
	wire   [31:0] mm_interconnect_0_parameter_sys_mapped_slave_writedata;         // mm_interconnect_0:Parameter_SYS_mapped_slave_writedata -> Parameter_SYS:mapped_slave_writedata
	wire    [0:0] mm_interconnect_0_parameter_sys_mapped_slave_burstcount;        // mm_interconnect_0:Parameter_SYS_mapped_slave_burstcount -> Parameter_SYS:mapped_slave_burstcount
	wire   [31:0] mm_interconnect_0_altpll_sys_pll_slave_readdata;                // altpll_sys:readdata -> mm_interconnect_0:altpll_sys_pll_slave_readdata
	wire    [1:0] mm_interconnect_0_altpll_sys_pll_slave_address;                 // mm_interconnect_0:altpll_sys_pll_slave_address -> altpll_sys:address
	wire          mm_interconnect_0_altpll_sys_pll_slave_read;                    // mm_interconnect_0:altpll_sys_pll_slave_read -> altpll_sys:read
	wire          mm_interconnect_0_altpll_sys_pll_slave_write;                   // mm_interconnect_0:altpll_sys_pll_slave_write -> altpll_sys:write
	wire   [31:0] mm_interconnect_0_altpll_sys_pll_slave_writedata;               // mm_interconnect_0:altpll_sys_pll_slave_writedata -> altpll_sys:writedata
	wire          mm_interconnect_0_program_memory_s1_chipselect;                 // mm_interconnect_0:Program_Memory_s1_chipselect -> Program_Memory:chipselect
	wire   [31:0] mm_interconnect_0_program_memory_s1_readdata;                   // Program_Memory:readdata -> mm_interconnect_0:Program_Memory_s1_readdata
	wire   [11:0] mm_interconnect_0_program_memory_s1_address;                    // mm_interconnect_0:Program_Memory_s1_address -> Program_Memory:address
	wire    [3:0] mm_interconnect_0_program_memory_s1_byteenable;                 // mm_interconnect_0:Program_Memory_s1_byteenable -> Program_Memory:byteenable
	wire          mm_interconnect_0_program_memory_s1_write;                      // mm_interconnect_0:Program_Memory_s1_write -> Program_Memory:write
	wire   [31:0] mm_interconnect_0_program_memory_s1_writedata;                  // mm_interconnect_0:Program_Memory_s1_writedata -> Program_Memory:writedata
	wire          mm_interconnect_0_program_memory_s1_clken;                      // mm_interconnect_0:Program_Memory_s1_clken -> Program_Memory:clken
	wire          mm_interconnect_0_data_memory_s1_chipselect;                    // mm_interconnect_0:Data_Memory_s1_chipselect -> Data_Memory:chipselect
	wire   [31:0] mm_interconnect_0_data_memory_s1_readdata;                      // Data_Memory:readdata -> mm_interconnect_0:Data_Memory_s1_readdata
	wire   [14:0] mm_interconnect_0_data_memory_s1_address;                       // mm_interconnect_0:Data_Memory_s1_address -> Data_Memory:address
	wire    [3:0] mm_interconnect_0_data_memory_s1_byteenable;                    // mm_interconnect_0:Data_Memory_s1_byteenable -> Data_Memory:byteenable
	wire          mm_interconnect_0_data_memory_s1_write;                         // mm_interconnect_0:Data_Memory_s1_write -> Data_Memory:write
	wire   [31:0] mm_interconnect_0_data_memory_s1_writedata;                     // mm_interconnect_0:Data_Memory_s1_writedata -> Data_Memory:writedata
	wire          mm_interconnect_0_data_memory_s1_clken;                         // mm_interconnect_0:Data_Memory_s1_clken -> Data_Memory:clken
	wire          irq_mapper_receiver0_irq;                                       // msgdma_0:csr_irq_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                       // external_bus_bridge:avalon_irq -> irq_mapper:receiver1_irq
	wire    [8:0] vic_0_irq_input_irq;                                            // irq_mapper:sender_irq -> vic_0:irq_input_irq
	wire          irq_mapper_receiver2_irq;                                       // irq_synchronizer:sender_irq -> irq_mapper:receiver2_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                                  // Parameter_SYS:parameter_loop_gpio_irq_irq -> irq_synchronizer:receiver_irq
	wire          irq_mapper_receiver3_irq;                                       // irq_synchronizer_001:sender_irq -> irq_mapper:receiver3_irq
	wire    [0:0] irq_synchronizer_001_receiver_irq;                              // TimerSYS_0:timer_0_irq_irq -> irq_synchronizer_001:receiver_irq
	wire          irq_mapper_receiver4_irq;                                       // irq_synchronizer_002:sender_irq -> irq_mapper:receiver4_irq
	wire    [0:0] irq_synchronizer_002_receiver_irq;                              // TimerSYS_0:timer_1_irq_irq -> irq_synchronizer_002:receiver_irq
	wire          rst_controller_reset_out_reset;                                 // rst_controller:reset_out -> [Data_Memory:reset, Parameter_SYS:slave_reset_reset, Pheriphals:slave_reset_reset, Program_Memory:reset, TimerSYS_0:slave_reset_reset, external_bus_bridge:reset, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, mm_interconnect_0:msgdma_0_reset_n_reset_bridge_in_reset_reset, msgdma_0:reset_n_reset_n, rst_translator:in_reset, vic_0:reset_reset]
	wire          rst_controller_reset_out_reset_req;                             // rst_controller:reset_req -> [Data_Memory:reset_req, Program_Memory:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_001_reset_out_reset;                             // rst_controller_001:reset_out -> [altpll_sys:reset, irq_synchronizer_001:receiver_reset, irq_synchronizer_002:receiver_reset, mm_interconnect_0:altpll_sys_inclk_interface_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_002_reset_out_reset;                             // rst_controller_002:reset_out -> [mm_interconnect_0:nios2_gen2_reset_reset_bridge_in_reset_reset, nios2_gen2:reset_n]
	wire          rst_controller_002_reset_out_reset_req;                         // rst_controller_002:reset_req -> nios2_gen2:reset_req
	wire          nios2_gen2_debug_reset_request_reset;                           // nios2_gen2:debug_reset_request -> rst_controller_002:reset_in1

	Mk8_Observer_CPU_Data_Memory data_memory (
		.clk        (cpu_clk_clk),                                 //   clk1.clk
		.address    (mm_interconnect_0_data_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_data_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_data_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_data_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_data_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_data_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_data_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),              // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),          //       .reset_req
		.freeze     (1'b0)                                         // (terminated)
	);

	Mk8_Observer_CPU_Parameter_SYS parameter_sys (
		.mapped_slave_waitrequest       (mm_interconnect_0_parameter_sys_mapped_slave_waitrequest),   //            mapped_slave.waitrequest
		.mapped_slave_readdata          (mm_interconnect_0_parameter_sys_mapped_slave_readdata),      //                        .readdata
		.mapped_slave_readdatavalid     (mm_interconnect_0_parameter_sys_mapped_slave_readdatavalid), //                        .readdatavalid
		.mapped_slave_burstcount        (mm_interconnect_0_parameter_sys_mapped_slave_burstcount),    //                        .burstcount
		.mapped_slave_writedata         (mm_interconnect_0_parameter_sys_mapped_slave_writedata),     //                        .writedata
		.mapped_slave_address           (mm_interconnect_0_parameter_sys_mapped_slave_address),       //                        .address
		.mapped_slave_write             (mm_interconnect_0_parameter_sys_mapped_slave_write),         //                        .write
		.mapped_slave_read              (mm_interconnect_0_parameter_sys_mapped_slave_read),          //                        .read
		.mapped_slave_byteenable        (mm_interconnect_0_parameter_sys_mapped_slave_byteenable),    //                        .byteenable
		.mapped_slave_debugaccess       (mm_interconnect_0_parameter_sys_mapped_slave_debugaccess),   //                        .debugaccess
		.parameter_clk_clk              (clk_clk),                                                    //           parameter_clk.clk
		.parameter_loop_gpio_in_port    (parameter_sys_parameter_loop_gpio_in_port),                  //     parameter_loop_gpio.in_port
		.parameter_loop_gpio_out_port   (parameter_sys_parameter_loop_gpio_out_port),                 //                        .out_port
		.parameter_loop_gpio_irq_irq    (irq_synchronizer_receiver_irq),                              // parameter_loop_gpio_irq.irq
		.parameter_reset_reset_n        (reset_reset_n),                                              //         parameter_reset.reset_n
		.parameter_rx_ram_s2_address    (parameter_sys_parameter_rx_ram_s2_address),                  //     parameter_rx_ram_s2.address
		.parameter_rx_ram_s2_chipselect (parameter_sys_parameter_rx_ram_s2_chipselect),               //                        .chipselect
		.parameter_rx_ram_s2_clken      (parameter_sys_parameter_rx_ram_s2_clken),                    //                        .clken
		.parameter_rx_ram_s2_write      (parameter_sys_parameter_rx_ram_s2_write),                    //                        .write
		.parameter_rx_ram_s2_readdata   (parameter_sys_parameter_rx_ram_s2_readdata),                 //                        .readdata
		.parameter_rx_ram_s2_writedata  (parameter_sys_parameter_rx_ram_s2_writedata),                //                        .writedata
		.parameter_rx_ram_s2_byteenable (parameter_sys_parameter_rx_ram_s2_byteenable),               //                        .byteenable
		.parameter_tx_ram_s2_address    (parameter_sys_parameter_tx_ram_s2_address),                  //     parameter_tx_ram_s2.address
		.parameter_tx_ram_s2_chipselect (parameter_sys_parameter_tx_ram_s2_chipselect),               //                        .chipselect
		.parameter_tx_ram_s2_clken      (parameter_sys_parameter_tx_ram_s2_clken),                    //                        .clken
		.parameter_tx_ram_s2_write      (parameter_sys_parameter_tx_ram_s2_write),                    //                        .write
		.parameter_tx_ram_s2_readdata   (parameter_sys_parameter_tx_ram_s2_readdata),                 //                        .readdata
		.parameter_tx_ram_s2_writedata  (parameter_sys_parameter_tx_ram_s2_writedata),                //                        .writedata
		.parameter_tx_ram_s2_byteenable (parameter_sys_parameter_tx_ram_s2_byteenable),               //                        .byteenable
		.pheriphal_clk_clk              (parameter_clk_1_clk),                                        //           pheriphal_clk.clk
		.pheriphal_reset_reset_n        (reset_parameter_reset_n),                                    //         pheriphal_reset.reset_n
		.reset_out_export               (parameter_sys_reset_out_export),                             //               reset_out.export
		.slave_clk_clk                  (cpu_clk_clk),                                                //               slave_clk.clk
		.slave_reset_reset              (rst_controller_reset_out_reset)                              //             slave_reset.reset
	);

	Mk8_Observer_CPU_Pheriphals pheriphals (
		.led_gpio_external_connection_export (pheriphals_led_gpio_external_connection_export),          // led_gpio_external_connection.export
		.mapped_slave_waitrequest            (mm_interconnect_0_pheriphals_mapped_slave_waitrequest),   //                 mapped_slave.waitrequest
		.mapped_slave_readdata               (mm_interconnect_0_pheriphals_mapped_slave_readdata),      //                             .readdata
		.mapped_slave_readdatavalid          (mm_interconnect_0_pheriphals_mapped_slave_readdatavalid), //                             .readdatavalid
		.mapped_slave_burstcount             (mm_interconnect_0_pheriphals_mapped_slave_burstcount),    //                             .burstcount
		.mapped_slave_writedata              (mm_interconnect_0_pheriphals_mapped_slave_writedata),     //                             .writedata
		.mapped_slave_address                (mm_interconnect_0_pheriphals_mapped_slave_address),       //                             .address
		.mapped_slave_write                  (mm_interconnect_0_pheriphals_mapped_slave_write),         //                             .write
		.mapped_slave_read                   (mm_interconnect_0_pheriphals_mapped_slave_read),          //                             .read
		.mapped_slave_byteenable             (mm_interconnect_0_pheriphals_mapped_slave_byteenable),    //                             .byteenable
		.mapped_slave_debugaccess            (mm_interconnect_0_pheriphals_mapped_slave_debugaccess),   //                             .debugaccess
		.pheriphal_clk_clk                   (clk_clk),                                                 //                pheriphal_clk.clk
		.pheriphal_reset_reset_n             (reset_reset_n),                                           //              pheriphal_reset.reset_n
		.slave_clk_clk                       (cpu_clk_clk),                                             //                    slave_clk.clk
		.slave_reset_reset                   (rst_controller_reset_out_reset),                          //                  slave_reset.reset
		.tp_gpio_external_connection_export  (pheriphals_tp_gpio_external_connection_export)            //  tp_gpio_external_connection.export
	);

	Mk8_Observer_CPU_Program_Memory program_memory (
		.clk        (cpu_clk_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_program_memory_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_program_memory_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_program_memory_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_program_memory_s1_write),      //       .write
		.readdata   (mm_interconnect_0_program_memory_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_program_memory_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_program_memory_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),                 // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),             //       .reset_req
		.freeze     (1'b0)                                            // (terminated)
	);

	Mk8_Observer_CPU_TimerSYS_0 timersys_0 (
		.mapped_slave_waitrequest   (mm_interconnect_0_timersys_0_mapped_slave_waitrequest),   //    mapped_slave.waitrequest
		.mapped_slave_readdata      (mm_interconnect_0_timersys_0_mapped_slave_readdata),      //                .readdata
		.mapped_slave_readdatavalid (mm_interconnect_0_timersys_0_mapped_slave_readdatavalid), //                .readdatavalid
		.mapped_slave_burstcount    (mm_interconnect_0_timersys_0_mapped_slave_burstcount),    //                .burstcount
		.mapped_slave_writedata     (mm_interconnect_0_timersys_0_mapped_slave_writedata),     //                .writedata
		.mapped_slave_address       (mm_interconnect_0_timersys_0_mapped_slave_address),       //                .address
		.mapped_slave_write         (mm_interconnect_0_timersys_0_mapped_slave_write),         //                .write
		.mapped_slave_read          (mm_interconnect_0_timersys_0_mapped_slave_read),          //                .read
		.mapped_slave_byteenable    (mm_interconnect_0_timersys_0_mapped_slave_byteenable),    //                .byteenable
		.mapped_slave_debugaccess   (mm_interconnect_0_timersys_0_mapped_slave_debugaccess),   //                .debugaccess
		.pheriphal_clk_clk          (clk_clk),                                                 //   pheriphal_clk.clk
		.pheriphal_reset_reset_n    (reset_reset_n),                                           // pheriphal_reset.reset_n
		.slave_clk_clk              (cpu_clk_clk),                                             //       slave_clk.clk
		.slave_reset_reset          (rst_controller_reset_out_reset),                          //     slave_reset.reset
		.timer_0_irq_irq            (irq_synchronizer_001_receiver_irq),                       //     timer_0_irq.irq
		.timer_1_irq_irq            (irq_synchronizer_002_receiver_irq)                        //     timer_1_irq.irq
	);

	Mk8_Observer_CPU_altpll_sys altpll_sys (
		.clk                (clk_clk),                                          //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),               // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_sys_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_sys_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_sys_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_sys_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_sys_pll_slave_writedata), //                      .writedata
		.c0                 (cpu_clk_clk),                                      //                    c0.clk
		.c1                 (clk_100m_clk),                                     //                    c1.clk
		.c2                 (clk_200m_clk),                                     //                    c2.clk
		.areset             (altpll_sys_areset_conduit_export),                 //        areset_conduit.export
		.locked             (altpll_sys_locked_conduit_export),                 //        locked_conduit.export
		.scandone           (),                                                 //           (terminated)
		.scandataout        (),                                                 //           (terminated)
		.c3                 (),                                                 //           (terminated)
		.c4                 (),                                                 //           (terminated)
		.phasedone          (),                                                 //           (terminated)
		.phasecounterselect (3'b000),                                           //           (terminated)
		.phaseupdown        (1'b0),                                             //           (terminated)
		.phasestep          (1'b0),                                             //           (terminated)
		.scanclk            (1'b0),                                             //           (terminated)
		.scanclkena         (1'b0),                                             //           (terminated)
		.scandata           (1'b0),                                             //           (terminated)
		.configupdate       (1'b0)                                              //           (terminated)
	);

	Mk8_Observer_CPU_external_bus_bridge external_bus_bridge (
		.clk                (cpu_clk_clk),                                                    //                clk.clk
		.reset              (rst_controller_reset_out_reset),                                 //              reset.reset
		.avalon_address     (mm_interconnect_0_external_bus_bridge_avalon_slave_address),     //       avalon_slave.address
		.avalon_byteenable  (mm_interconnect_0_external_bus_bridge_avalon_slave_byteenable),  //                   .byteenable
		.avalon_chipselect  (mm_interconnect_0_external_bus_bridge_avalon_slave_chipselect),  //                   .chipselect
		.avalon_read        (mm_interconnect_0_external_bus_bridge_avalon_slave_read),        //                   .read
		.avalon_write       (mm_interconnect_0_external_bus_bridge_avalon_slave_write),       //                   .write
		.avalon_writedata   (mm_interconnect_0_external_bus_bridge_avalon_slave_writedata),   //                   .writedata
		.avalon_readdata    (mm_interconnect_0_external_bus_bridge_avalon_slave_readdata),    //                   .readdata
		.avalon_waitrequest (mm_interconnect_0_external_bus_bridge_avalon_slave_waitrequest), //                   .waitrequest
		.avalon_irq         (irq_mapper_receiver1_irq),                                       //          interrupt.irq
		.acknowledge        (external_bus_bridge_external_interface_acknowledge),             // external_interface.export
		.irq                (external_bus_bridge_external_interface_irq),                     //                   .export
		.address            (external_bus_bridge_external_interface_address),                 //                   .export
		.bus_enable         (external_bus_bridge_external_interface_bus_enable),              //                   .export
		.byte_enable        (external_bus_bridge_external_interface_byte_enable),             //                   .export
		.rw                 (external_bus_bridge_external_interface_rw),                      //                   .export
		.write_data         (external_bus_bridge_external_interface_write_data),              //                   .export
		.read_data          (external_bus_bridge_external_interface_read_data)                //                   .export
	);

	Mk8_Observer_CPU_msgdma_0 msgdma_0 (
		.mm_read_address              (msgdma_0_mm_read_address),                                //          mm_read.address
		.mm_read_read                 (msgdma_0_mm_read_read),                                   //                 .read
		.mm_read_byteenable           (msgdma_0_mm_read_byteenable),                             //                 .byteenable
		.mm_read_readdata             (msgdma_0_mm_read_readdata),                               //                 .readdata
		.mm_read_waitrequest          (msgdma_0_mm_read_waitrequest),                            //                 .waitrequest
		.mm_read_readdatavalid        (msgdma_0_mm_read_readdatavalid),                          //                 .readdatavalid
		.mm_write_address             (msgdma_0_mm_write_address),                               //         mm_write.address
		.mm_write_write               (msgdma_0_mm_write_write),                                 //                 .write
		.mm_write_byteenable          (msgdma_0_mm_write_byteenable),                            //                 .byteenable
		.mm_write_writedata           (msgdma_0_mm_write_writedata),                             //                 .writedata
		.mm_write_waitrequest         (msgdma_0_mm_write_waitrequest),                           //                 .waitrequest
		.clock_clk                    (cpu_clk_clk),                                             //            clock.clk
		.reset_n_reset_n              (~rst_controller_reset_out_reset),                         //          reset_n.reset_n
		.csr_writedata                (mm_interconnect_0_msgdma_0_csr_writedata),                //              csr.writedata
		.csr_write                    (mm_interconnect_0_msgdma_0_csr_write),                    //                 .write
		.csr_byteenable               (mm_interconnect_0_msgdma_0_csr_byteenable),               //                 .byteenable
		.csr_readdata                 (mm_interconnect_0_msgdma_0_csr_readdata),                 //                 .readdata
		.csr_read                     (mm_interconnect_0_msgdma_0_csr_read),                     //                 .read
		.csr_address                  (mm_interconnect_0_msgdma_0_csr_address),                  //                 .address
		.descriptor_slave_write       (mm_interconnect_0_msgdma_0_descriptor_slave_write),       // descriptor_slave.write
		.descriptor_slave_waitrequest (mm_interconnect_0_msgdma_0_descriptor_slave_waitrequest), //                 .waitrequest
		.descriptor_slave_writedata   (mm_interconnect_0_msgdma_0_descriptor_slave_writedata),   //                 .writedata
		.descriptor_slave_byteenable  (mm_interconnect_0_msgdma_0_descriptor_slave_byteenable),  //                 .byteenable
		.csr_irq_irq                  (irq_mapper_receiver0_irq)                                 //          csr_irq.irq
	);

	Mk8_Observer_CPU_nios2_gen2 nios2_gen2 (
		.clk                                 (cpu_clk_clk),                                              //                       clk.clk
		.reset_n                             (~rst_controller_002_reset_out_reset),                      //                     reset.reset_n
		.reset_req                           (rst_controller_002_reset_out_reset_req),                   //                          .reset_req
		.d_address                           (nios2_gen2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (nios2_gen2_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (nios2_gen2_instruction_master_readdatavalid),              //                          .readdatavalid
		.eic_port_valid                      (vic_0_interrupt_controller_out_valid),                     //   interrupt_controller_in.valid
		.eic_port_data                       (vic_0_interrupt_controller_out_data),                      //                          .data
		.debug_reset_request                 (nios2_gen2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                          // custom_instruction_master.readra
	);

	Mk8_Observer_CPU_vic_0 vic_0 (
		.clk_clk                        (cpu_clk_clk),                                  //                      clk.clk
		.reset_reset                    (rst_controller_reset_out_reset),               //                    reset.reset
		.irq_input_irq                  (vic_0_irq_input_irq),                          //                irq_input.irq
		.csr_access_read                (mm_interconnect_0_vic_0_csr_access_read),      //               csr_access.read
		.csr_access_write               (mm_interconnect_0_vic_0_csr_access_write),     //                         .write
		.csr_access_address             (mm_interconnect_0_vic_0_csr_access_address),   //                         .address
		.csr_access_writedata           (mm_interconnect_0_vic_0_csr_access_writedata), //                         .writedata
		.csr_access_readdata            (mm_interconnect_0_vic_0_csr_access_readdata),  //                         .readdata
		.interrupt_controller_out_valid (vic_0_interrupt_controller_out_valid),         // interrupt_controller_out.valid
		.interrupt_controller_out_data  (vic_0_interrupt_controller_out_data)           //                         .data
	);

	Mk8_Observer_CPU_mm_interconnect_0 mm_interconnect_0 (
		.altpll_sys_c0_clk                                            (cpu_clk_clk),                                                    //                                          altpll_sys_c0.clk
		.clk_50_clk_clk                                               (clk_clk),                                                        //                                             clk_50_clk.clk
		.altpll_sys_inclk_interface_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                             // altpll_sys_inclk_interface_reset_reset_bridge_in_reset.reset
		.msgdma_0_reset_n_reset_bridge_in_reset_reset                 (rst_controller_reset_out_reset),                                 //                 msgdma_0_reset_n_reset_bridge_in_reset.reset
		.nios2_gen2_reset_reset_bridge_in_reset_reset                 (rst_controller_002_reset_out_reset),                             //                 nios2_gen2_reset_reset_bridge_in_reset.reset
		.msgdma_0_mm_read_address                                     (msgdma_0_mm_read_address),                                       //                                       msgdma_0_mm_read.address
		.msgdma_0_mm_read_waitrequest                                 (msgdma_0_mm_read_waitrequest),                                   //                                                       .waitrequest
		.msgdma_0_mm_read_byteenable                                  (msgdma_0_mm_read_byteenable),                                    //                                                       .byteenable
		.msgdma_0_mm_read_read                                        (msgdma_0_mm_read_read),                                          //                                                       .read
		.msgdma_0_mm_read_readdata                                    (msgdma_0_mm_read_readdata),                                      //                                                       .readdata
		.msgdma_0_mm_read_readdatavalid                               (msgdma_0_mm_read_readdatavalid),                                 //                                                       .readdatavalid
		.msgdma_0_mm_write_address                                    (msgdma_0_mm_write_address),                                      //                                      msgdma_0_mm_write.address
		.msgdma_0_mm_write_waitrequest                                (msgdma_0_mm_write_waitrequest),                                  //                                                       .waitrequest
		.msgdma_0_mm_write_byteenable                                 (msgdma_0_mm_write_byteenable),                                   //                                                       .byteenable
		.msgdma_0_mm_write_write                                      (msgdma_0_mm_write_write),                                        //                                                       .write
		.msgdma_0_mm_write_writedata                                  (msgdma_0_mm_write_writedata),                                    //                                                       .writedata
		.nios2_gen2_data_master_address                               (nios2_gen2_data_master_address),                                 //                                 nios2_gen2_data_master.address
		.nios2_gen2_data_master_waitrequest                           (nios2_gen2_data_master_waitrequest),                             //                                                       .waitrequest
		.nios2_gen2_data_master_byteenable                            (nios2_gen2_data_master_byteenable),                              //                                                       .byteenable
		.nios2_gen2_data_master_read                                  (nios2_gen2_data_master_read),                                    //                                                       .read
		.nios2_gen2_data_master_readdata                              (nios2_gen2_data_master_readdata),                                //                                                       .readdata
		.nios2_gen2_data_master_readdatavalid                         (nios2_gen2_data_master_readdatavalid),                           //                                                       .readdatavalid
		.nios2_gen2_data_master_write                                 (nios2_gen2_data_master_write),                                   //                                                       .write
		.nios2_gen2_data_master_writedata                             (nios2_gen2_data_master_writedata),                               //                                                       .writedata
		.nios2_gen2_data_master_debugaccess                           (nios2_gen2_data_master_debugaccess),                             //                                                       .debugaccess
		.nios2_gen2_instruction_master_address                        (nios2_gen2_instruction_master_address),                          //                          nios2_gen2_instruction_master.address
		.nios2_gen2_instruction_master_waitrequest                    (nios2_gen2_instruction_master_waitrequest),                      //                                                       .waitrequest
		.nios2_gen2_instruction_master_read                           (nios2_gen2_instruction_master_read),                             //                                                       .read
		.nios2_gen2_instruction_master_readdata                       (nios2_gen2_instruction_master_readdata),                         //                                                       .readdata
		.nios2_gen2_instruction_master_readdatavalid                  (nios2_gen2_instruction_master_readdatavalid),                    //                                                       .readdatavalid
		.altpll_sys_pll_slave_address                                 (mm_interconnect_0_altpll_sys_pll_slave_address),                 //                                   altpll_sys_pll_slave.address
		.altpll_sys_pll_slave_write                                   (mm_interconnect_0_altpll_sys_pll_slave_write),                   //                                                       .write
		.altpll_sys_pll_slave_read                                    (mm_interconnect_0_altpll_sys_pll_slave_read),                    //                                                       .read
		.altpll_sys_pll_slave_readdata                                (mm_interconnect_0_altpll_sys_pll_slave_readdata),                //                                                       .readdata
		.altpll_sys_pll_slave_writedata                               (mm_interconnect_0_altpll_sys_pll_slave_writedata),               //                                                       .writedata
		.Data_Memory_s1_address                                       (mm_interconnect_0_data_memory_s1_address),                       //                                         Data_Memory_s1.address
		.Data_Memory_s1_write                                         (mm_interconnect_0_data_memory_s1_write),                         //                                                       .write
		.Data_Memory_s1_readdata                                      (mm_interconnect_0_data_memory_s1_readdata),                      //                                                       .readdata
		.Data_Memory_s1_writedata                                     (mm_interconnect_0_data_memory_s1_writedata),                     //                                                       .writedata
		.Data_Memory_s1_byteenable                                    (mm_interconnect_0_data_memory_s1_byteenable),                    //                                                       .byteenable
		.Data_Memory_s1_chipselect                                    (mm_interconnect_0_data_memory_s1_chipselect),                    //                                                       .chipselect
		.Data_Memory_s1_clken                                         (mm_interconnect_0_data_memory_s1_clken),                         //                                                       .clken
		.external_bus_bridge_avalon_slave_address                     (mm_interconnect_0_external_bus_bridge_avalon_slave_address),     //                       external_bus_bridge_avalon_slave.address
		.external_bus_bridge_avalon_slave_write                       (mm_interconnect_0_external_bus_bridge_avalon_slave_write),       //                                                       .write
		.external_bus_bridge_avalon_slave_read                        (mm_interconnect_0_external_bus_bridge_avalon_slave_read),        //                                                       .read
		.external_bus_bridge_avalon_slave_readdata                    (mm_interconnect_0_external_bus_bridge_avalon_slave_readdata),    //                                                       .readdata
		.external_bus_bridge_avalon_slave_writedata                   (mm_interconnect_0_external_bus_bridge_avalon_slave_writedata),   //                                                       .writedata
		.external_bus_bridge_avalon_slave_byteenable                  (mm_interconnect_0_external_bus_bridge_avalon_slave_byteenable),  //                                                       .byteenable
		.external_bus_bridge_avalon_slave_waitrequest                 (mm_interconnect_0_external_bus_bridge_avalon_slave_waitrequest), //                                                       .waitrequest
		.external_bus_bridge_avalon_slave_chipselect                  (mm_interconnect_0_external_bus_bridge_avalon_slave_chipselect),  //                                                       .chipselect
		.msgdma_0_csr_address                                         (mm_interconnect_0_msgdma_0_csr_address),                         //                                           msgdma_0_csr.address
		.msgdma_0_csr_write                                           (mm_interconnect_0_msgdma_0_csr_write),                           //                                                       .write
		.msgdma_0_csr_read                                            (mm_interconnect_0_msgdma_0_csr_read),                            //                                                       .read
		.msgdma_0_csr_readdata                                        (mm_interconnect_0_msgdma_0_csr_readdata),                        //                                                       .readdata
		.msgdma_0_csr_writedata                                       (mm_interconnect_0_msgdma_0_csr_writedata),                       //                                                       .writedata
		.msgdma_0_csr_byteenable                                      (mm_interconnect_0_msgdma_0_csr_byteenable),                      //                                                       .byteenable
		.msgdma_0_descriptor_slave_write                              (mm_interconnect_0_msgdma_0_descriptor_slave_write),              //                              msgdma_0_descriptor_slave.write
		.msgdma_0_descriptor_slave_writedata                          (mm_interconnect_0_msgdma_0_descriptor_slave_writedata),          //                                                       .writedata
		.msgdma_0_descriptor_slave_byteenable                         (mm_interconnect_0_msgdma_0_descriptor_slave_byteenable),         //                                                       .byteenable
		.msgdma_0_descriptor_slave_waitrequest                        (mm_interconnect_0_msgdma_0_descriptor_slave_waitrequest),        //                                                       .waitrequest
		.nios2_gen2_debug_mem_slave_address                           (mm_interconnect_0_nios2_gen2_debug_mem_slave_address),           //                             nios2_gen2_debug_mem_slave.address
		.nios2_gen2_debug_mem_slave_write                             (mm_interconnect_0_nios2_gen2_debug_mem_slave_write),             //                                                       .write
		.nios2_gen2_debug_mem_slave_read                              (mm_interconnect_0_nios2_gen2_debug_mem_slave_read),              //                                                       .read
		.nios2_gen2_debug_mem_slave_readdata                          (mm_interconnect_0_nios2_gen2_debug_mem_slave_readdata),          //                                                       .readdata
		.nios2_gen2_debug_mem_slave_writedata                         (mm_interconnect_0_nios2_gen2_debug_mem_slave_writedata),         //                                                       .writedata
		.nios2_gen2_debug_mem_slave_byteenable                        (mm_interconnect_0_nios2_gen2_debug_mem_slave_byteenable),        //                                                       .byteenable
		.nios2_gen2_debug_mem_slave_waitrequest                       (mm_interconnect_0_nios2_gen2_debug_mem_slave_waitrequest),       //                                                       .waitrequest
		.nios2_gen2_debug_mem_slave_debugaccess                       (mm_interconnect_0_nios2_gen2_debug_mem_slave_debugaccess),       //                                                       .debugaccess
		.Parameter_SYS_mapped_slave_address                           (mm_interconnect_0_parameter_sys_mapped_slave_address),           //                             Parameter_SYS_mapped_slave.address
		.Parameter_SYS_mapped_slave_write                             (mm_interconnect_0_parameter_sys_mapped_slave_write),             //                                                       .write
		.Parameter_SYS_mapped_slave_read                              (mm_interconnect_0_parameter_sys_mapped_slave_read),              //                                                       .read
		.Parameter_SYS_mapped_slave_readdata                          (mm_interconnect_0_parameter_sys_mapped_slave_readdata),          //                                                       .readdata
		.Parameter_SYS_mapped_slave_writedata                         (mm_interconnect_0_parameter_sys_mapped_slave_writedata),         //                                                       .writedata
		.Parameter_SYS_mapped_slave_burstcount                        (mm_interconnect_0_parameter_sys_mapped_slave_burstcount),        //                                                       .burstcount
		.Parameter_SYS_mapped_slave_byteenable                        (mm_interconnect_0_parameter_sys_mapped_slave_byteenable),        //                                                       .byteenable
		.Parameter_SYS_mapped_slave_readdatavalid                     (mm_interconnect_0_parameter_sys_mapped_slave_readdatavalid),     //                                                       .readdatavalid
		.Parameter_SYS_mapped_slave_waitrequest                       (mm_interconnect_0_parameter_sys_mapped_slave_waitrequest),       //                                                       .waitrequest
		.Parameter_SYS_mapped_slave_debugaccess                       (mm_interconnect_0_parameter_sys_mapped_slave_debugaccess),       //                                                       .debugaccess
		.Pheriphals_mapped_slave_address                              (mm_interconnect_0_pheriphals_mapped_slave_address),              //                                Pheriphals_mapped_slave.address
		.Pheriphals_mapped_slave_write                                (mm_interconnect_0_pheriphals_mapped_slave_write),                //                                                       .write
		.Pheriphals_mapped_slave_read                                 (mm_interconnect_0_pheriphals_mapped_slave_read),                 //                                                       .read
		.Pheriphals_mapped_slave_readdata                             (mm_interconnect_0_pheriphals_mapped_slave_readdata),             //                                                       .readdata
		.Pheriphals_mapped_slave_writedata                            (mm_interconnect_0_pheriphals_mapped_slave_writedata),            //                                                       .writedata
		.Pheriphals_mapped_slave_burstcount                           (mm_interconnect_0_pheriphals_mapped_slave_burstcount),           //                                                       .burstcount
		.Pheriphals_mapped_slave_byteenable                           (mm_interconnect_0_pheriphals_mapped_slave_byteenable),           //                                                       .byteenable
		.Pheriphals_mapped_slave_readdatavalid                        (mm_interconnect_0_pheriphals_mapped_slave_readdatavalid),        //                                                       .readdatavalid
		.Pheriphals_mapped_slave_waitrequest                          (mm_interconnect_0_pheriphals_mapped_slave_waitrequest),          //                                                       .waitrequest
		.Pheriphals_mapped_slave_debugaccess                          (mm_interconnect_0_pheriphals_mapped_slave_debugaccess),          //                                                       .debugaccess
		.Program_Memory_s1_address                                    (mm_interconnect_0_program_memory_s1_address),                    //                                      Program_Memory_s1.address
		.Program_Memory_s1_write                                      (mm_interconnect_0_program_memory_s1_write),                      //                                                       .write
		.Program_Memory_s1_readdata                                   (mm_interconnect_0_program_memory_s1_readdata),                   //                                                       .readdata
		.Program_Memory_s1_writedata                                  (mm_interconnect_0_program_memory_s1_writedata),                  //                                                       .writedata
		.Program_Memory_s1_byteenable                                 (mm_interconnect_0_program_memory_s1_byteenable),                 //                                                       .byteenable
		.Program_Memory_s1_chipselect                                 (mm_interconnect_0_program_memory_s1_chipselect),                 //                                                       .chipselect
		.Program_Memory_s1_clken                                      (mm_interconnect_0_program_memory_s1_clken),                      //                                                       .clken
		.TimerSYS_0_mapped_slave_address                              (mm_interconnect_0_timersys_0_mapped_slave_address),              //                                TimerSYS_0_mapped_slave.address
		.TimerSYS_0_mapped_slave_write                                (mm_interconnect_0_timersys_0_mapped_slave_write),                //                                                       .write
		.TimerSYS_0_mapped_slave_read                                 (mm_interconnect_0_timersys_0_mapped_slave_read),                 //                                                       .read
		.TimerSYS_0_mapped_slave_readdata                             (mm_interconnect_0_timersys_0_mapped_slave_readdata),             //                                                       .readdata
		.TimerSYS_0_mapped_slave_writedata                            (mm_interconnect_0_timersys_0_mapped_slave_writedata),            //                                                       .writedata
		.TimerSYS_0_mapped_slave_burstcount                           (mm_interconnect_0_timersys_0_mapped_slave_burstcount),           //                                                       .burstcount
		.TimerSYS_0_mapped_slave_byteenable                           (mm_interconnect_0_timersys_0_mapped_slave_byteenable),           //                                                       .byteenable
		.TimerSYS_0_mapped_slave_readdatavalid                        (mm_interconnect_0_timersys_0_mapped_slave_readdatavalid),        //                                                       .readdatavalid
		.TimerSYS_0_mapped_slave_waitrequest                          (mm_interconnect_0_timersys_0_mapped_slave_waitrequest),          //                                                       .waitrequest
		.TimerSYS_0_mapped_slave_debugaccess                          (mm_interconnect_0_timersys_0_mapped_slave_debugaccess),          //                                                       .debugaccess
		.vic_0_csr_access_address                                     (mm_interconnect_0_vic_0_csr_access_address),                     //                                       vic_0_csr_access.address
		.vic_0_csr_access_write                                       (mm_interconnect_0_vic_0_csr_access_write),                       //                                                       .write
		.vic_0_csr_access_read                                        (mm_interconnect_0_vic_0_csr_access_read),                        //                                                       .read
		.vic_0_csr_access_readdata                                    (mm_interconnect_0_vic_0_csr_access_readdata),                    //                                                       .readdata
		.vic_0_csr_access_writedata                                   (mm_interconnect_0_vic_0_csr_access_writedata)                    //                                                       .writedata
	);

	Mk8_Observer_CPU_irq_mapper irq_mapper (
		.clk           (cpu_clk_clk),                    //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),       // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),       // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),       // receiver4.irq
		.sender_irq    (vic_0_irq_input_irq)             //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (cpu_clk_clk),                    //       receiver_clk.clk
		.sender_clk     (cpu_clk_clk),                    //         sender_clk.clk
		.receiver_reset (),                               // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)        //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (cpu_clk_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (cpu_clk_clk),                        //         sender_clk.clk
		.receiver_reset (rst_controller_001_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_reset_out_reset),     //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (cpu_clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_debug_reset_request_reset),   // reset_in1.reset
		.clk            (cpu_clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
