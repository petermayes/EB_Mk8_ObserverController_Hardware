// Pararameter_Comms_SYS.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module Pararameter_Comms_SYS (
		output wire        mapped_slave_waitrequest,       //            mapped_slave.waitrequest
		output wire [31:0] mapped_slave_readdata,          //                        .readdata
		output wire        mapped_slave_readdatavalid,     //                        .readdatavalid
		input  wire [0:0]  mapped_slave_burstcount,        //                        .burstcount
		input  wire [31:0] mapped_slave_writedata,         //                        .writedata
		input  wire [14:0] mapped_slave_address,           //                        .address
		input  wire        mapped_slave_write,             //                        .write
		input  wire        mapped_slave_read,              //                        .read
		input  wire [3:0]  mapped_slave_byteenable,        //                        .byteenable
		input  wire        mapped_slave_debugaccess,       //                        .debugaccess
		input  wire        parameter_clk_clk,              //           parameter_clk.clk
		input  wire        parameter_loop_gpio_in_port,    //     parameter_loop_gpio.in_port
		output wire        parameter_loop_gpio_out_port,   //                        .out_port
		output wire        parameter_loop_gpio_irq_irq,    // parameter_loop_gpio_irq.irq
		input  wire        parameter_reset_reset_n,        //         parameter_reset.reset_n
		input  wire [10:0] parameter_rx_ram_s2_address,    //     parameter_rx_ram_s2.address
		input  wire        parameter_rx_ram_s2_chipselect, //                        .chipselect
		input  wire        parameter_rx_ram_s2_clken,      //                        .clken
		input  wire        parameter_rx_ram_s2_write,      //                        .write
		output wire [31:0] parameter_rx_ram_s2_readdata,   //                        .readdata
		input  wire [31:0] parameter_rx_ram_s2_writedata,  //                        .writedata
		input  wire [3:0]  parameter_rx_ram_s2_byteenable, //                        .byteenable
		input  wire [10:0] parameter_tx_ram_s2_address,    //     parameter_tx_ram_s2.address
		input  wire        parameter_tx_ram_s2_chipselect, //                        .chipselect
		input  wire        parameter_tx_ram_s2_clken,      //                        .clken
		input  wire        parameter_tx_ram_s2_write,      //                        .write
		output wire [31:0] parameter_tx_ram_s2_readdata,   //                        .readdata
		input  wire [31:0] parameter_tx_ram_s2_writedata,  //                        .writedata
		input  wire [3:0]  parameter_tx_ram_s2_byteenable, //                        .byteenable
		input  wire        pheriphal_clk_clk,              //           pheriphal_clk.clk
		input  wire        pheriphal_reset_reset_n,        //         pheriphal_reset.reset_n
		output wire        reset_out_export,               //               reset_out.export
		input  wire        slave_clk_clk,                  //               slave_clk.clk
		input  wire        slave_reset_reset               //             slave_reset.reset
	);

	wire         mm_clock_crossing_bridge_0_m0_waitrequest;        // mm_interconnect_0:mm_clock_crossing_bridge_0_m0_waitrequest -> mm_clock_crossing_bridge_0:m0_waitrequest
	wire  [31:0] mm_clock_crossing_bridge_0_m0_readdata;           // mm_interconnect_0:mm_clock_crossing_bridge_0_m0_readdata -> mm_clock_crossing_bridge_0:m0_readdata
	wire         mm_clock_crossing_bridge_0_m0_debugaccess;        // mm_clock_crossing_bridge_0:m0_debugaccess -> mm_interconnect_0:mm_clock_crossing_bridge_0_m0_debugaccess
	wire  [14:0] mm_clock_crossing_bridge_0_m0_address;            // mm_clock_crossing_bridge_0:m0_address -> mm_interconnect_0:mm_clock_crossing_bridge_0_m0_address
	wire         mm_clock_crossing_bridge_0_m0_read;               // mm_clock_crossing_bridge_0:m0_read -> mm_interconnect_0:mm_clock_crossing_bridge_0_m0_read
	wire   [3:0] mm_clock_crossing_bridge_0_m0_byteenable;         // mm_clock_crossing_bridge_0:m0_byteenable -> mm_interconnect_0:mm_clock_crossing_bridge_0_m0_byteenable
	wire         mm_clock_crossing_bridge_0_m0_readdatavalid;      // mm_interconnect_0:mm_clock_crossing_bridge_0_m0_readdatavalid -> mm_clock_crossing_bridge_0:m0_readdatavalid
	wire  [31:0] mm_clock_crossing_bridge_0_m0_writedata;          // mm_clock_crossing_bridge_0:m0_writedata -> mm_interconnect_0:mm_clock_crossing_bridge_0_m0_writedata
	wire         mm_clock_crossing_bridge_0_m0_write;              // mm_clock_crossing_bridge_0:m0_write -> mm_interconnect_0:mm_clock_crossing_bridge_0_m0_write
	wire   [0:0] mm_clock_crossing_bridge_0_m0_burstcount;         // mm_clock_crossing_bridge_0:m0_burstcount -> mm_interconnect_0:mm_clock_crossing_bridge_0_m0_burstcount
	wire         mm_interconnect_0_parameter_gpio_s1_chipselect;   // mm_interconnect_0:Parameter_GPIO_s1_chipselect -> Parameter_GPIO:chipselect
	wire  [31:0] mm_interconnect_0_parameter_gpio_s1_readdata;     // Parameter_GPIO:readdata -> mm_interconnect_0:Parameter_GPIO_s1_readdata
	wire   [2:0] mm_interconnect_0_parameter_gpio_s1_address;      // mm_interconnect_0:Parameter_GPIO_s1_address -> Parameter_GPIO:address
	wire         mm_interconnect_0_parameter_gpio_s1_write;        // mm_interconnect_0:Parameter_GPIO_s1_write -> Parameter_GPIO:write_n
	wire  [31:0] mm_interconnect_0_parameter_gpio_s1_writedata;    // mm_interconnect_0:Parameter_GPIO_s1_writedata -> Parameter_GPIO:writedata
	wire         mm_interconnect_0_parameter_rx_ram_s1_chipselect; // mm_interconnect_0:Parameter_RX_RAM_s1_chipselect -> Parameter_RX_RAM:chipselect
	wire  [31:0] mm_interconnect_0_parameter_rx_ram_s1_readdata;   // Parameter_RX_RAM:readdata -> mm_interconnect_0:Parameter_RX_RAM_s1_readdata
	wire  [10:0] mm_interconnect_0_parameter_rx_ram_s1_address;    // mm_interconnect_0:Parameter_RX_RAM_s1_address -> Parameter_RX_RAM:address
	wire   [3:0] mm_interconnect_0_parameter_rx_ram_s1_byteenable; // mm_interconnect_0:Parameter_RX_RAM_s1_byteenable -> Parameter_RX_RAM:byteenable
	wire         mm_interconnect_0_parameter_rx_ram_s1_write;      // mm_interconnect_0:Parameter_RX_RAM_s1_write -> Parameter_RX_RAM:write
	wire  [31:0] mm_interconnect_0_parameter_rx_ram_s1_writedata;  // mm_interconnect_0:Parameter_RX_RAM_s1_writedata -> Parameter_RX_RAM:writedata
	wire         mm_interconnect_0_parameter_rx_ram_s1_clken;      // mm_interconnect_0:Parameter_RX_RAM_s1_clken -> Parameter_RX_RAM:clken
	wire         mm_interconnect_0_reset_s1_chipselect;            // mm_interconnect_0:Reset_s1_chipselect -> Reset:chipselect
	wire  [31:0] mm_interconnect_0_reset_s1_readdata;              // Reset:readdata -> mm_interconnect_0:Reset_s1_readdata
	wire   [2:0] mm_interconnect_0_reset_s1_address;               // mm_interconnect_0:Reset_s1_address -> Reset:address
	wire         mm_interconnect_0_reset_s1_write;                 // mm_interconnect_0:Reset_s1_write -> Reset:write_n
	wire  [31:0] mm_interconnect_0_reset_s1_writedata;             // mm_interconnect_0:Reset_s1_writedata -> Reset:writedata
	wire         mm_interconnect_0_parameter_tx_ram_s1_chipselect; // mm_interconnect_0:Parameter_TX_RAM_s1_chipselect -> Parameter_TX_RAM:chipselect
	wire  [31:0] mm_interconnect_0_parameter_tx_ram_s1_readdata;   // Parameter_TX_RAM:readdata -> mm_interconnect_0:Parameter_TX_RAM_s1_readdata
	wire  [10:0] mm_interconnect_0_parameter_tx_ram_s1_address;    // mm_interconnect_0:Parameter_TX_RAM_s1_address -> Parameter_TX_RAM:address
	wire   [3:0] mm_interconnect_0_parameter_tx_ram_s1_byteenable; // mm_interconnect_0:Parameter_TX_RAM_s1_byteenable -> Parameter_TX_RAM:byteenable
	wire         mm_interconnect_0_parameter_tx_ram_s1_write;      // mm_interconnect_0:Parameter_TX_RAM_s1_write -> Parameter_TX_RAM:write
	wire  [31:0] mm_interconnect_0_parameter_tx_ram_s1_writedata;  // mm_interconnect_0:Parameter_TX_RAM_s1_writedata -> Parameter_TX_RAM:writedata
	wire         mm_interconnect_0_parameter_tx_ram_s1_clken;      // mm_interconnect_0:Parameter_TX_RAM_s1_clken -> Parameter_TX_RAM:clken
	wire         rst_controller_reset_out_reset;                   // rst_controller:reset_out -> [Parameter_GPIO:reset_n, Parameter_RX_RAM:reset, Parameter_TX_RAM:reset, Reset:reset_n, mm_clock_crossing_bridge_0:m0_reset, mm_interconnect_0:mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;               // rst_controller:reset_req -> [Parameter_RX_RAM:reset_req, Parameter_TX_RAM:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_001_reset_out_reset;               // rst_controller_001:reset_out -> [Parameter_RX_RAM:reset2, Parameter_TX_RAM:reset2]
	wire         rst_controller_001_reset_out_reset_req;           // rst_controller_001:reset_req -> [Parameter_RX_RAM:reset_req2, Parameter_TX_RAM:reset_req2]

	Pararameter_Comms_SYS_Parameter_GPIO parameter_gpio (
		.clk        (pheriphal_clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                //               reset.reset_n
		.address    (mm_interconnect_0_parameter_gpio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_parameter_gpio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_parameter_gpio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_parameter_gpio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_parameter_gpio_s1_readdata),   //                    .readdata
		.in_port    (parameter_loop_gpio_in_port),                    // external_connection.export
		.out_port   (parameter_loop_gpio_out_port),                   //                    .export
		.irq        (parameter_loop_gpio_irq_irq)                     //                 irq.irq
	);

	Pararameter_Comms_SYS_Parameter_RX_RAM parameter_rx_ram (
		.clk         (pheriphal_clk_clk),                                //   clk1.clk
		.address     (mm_interconnect_0_parameter_rx_ram_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_parameter_rx_ram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_parameter_rx_ram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_parameter_rx_ram_s1_write),      //       .write
		.readdata    (mm_interconnect_0_parameter_rx_ram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_parameter_rx_ram_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_parameter_rx_ram_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),               //       .reset_req
		.address2    (parameter_rx_ram_s2_address),                      //     s2.address
		.chipselect2 (parameter_rx_ram_s2_chipselect),                   //       .chipselect
		.clken2      (parameter_rx_ram_s2_clken),                        //       .clken
		.write2      (parameter_rx_ram_s2_write),                        //       .write
		.readdata2   (parameter_rx_ram_s2_readdata),                     //       .readdata
		.writedata2  (parameter_rx_ram_s2_writedata),                    //       .writedata
		.byteenable2 (parameter_rx_ram_s2_byteenable),                   //       .byteenable
		.clk2        (parameter_clk_clk),                                //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),               // reset2.reset
		.reset_req2  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze      (1'b0)                                              // (terminated)
	);

	Pararameter_Comms_SYS_Parameter_TX_RAM parameter_tx_ram (
		.clk         (pheriphal_clk_clk),                                //   clk1.clk
		.address     (mm_interconnect_0_parameter_tx_ram_s1_address),    //     s1.address
		.clken       (mm_interconnect_0_parameter_tx_ram_s1_clken),      //       .clken
		.chipselect  (mm_interconnect_0_parameter_tx_ram_s1_chipselect), //       .chipselect
		.write       (mm_interconnect_0_parameter_tx_ram_s1_write),      //       .write
		.readdata    (mm_interconnect_0_parameter_tx_ram_s1_readdata),   //       .readdata
		.writedata   (mm_interconnect_0_parameter_tx_ram_s1_writedata),  //       .writedata
		.byteenable  (mm_interconnect_0_parameter_tx_ram_s1_byteenable), //       .byteenable
		.reset       (rst_controller_reset_out_reset),                   // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),               //       .reset_req
		.address2    (parameter_tx_ram_s2_address),                      //     s2.address
		.chipselect2 (parameter_tx_ram_s2_chipselect),                   //       .chipselect
		.clken2      (parameter_tx_ram_s2_clken),                        //       .clken
		.write2      (parameter_tx_ram_s2_write),                        //       .write
		.readdata2   (parameter_tx_ram_s2_readdata),                     //       .readdata
		.writedata2  (parameter_tx_ram_s2_writedata),                    //       .writedata
		.byteenable2 (parameter_tx_ram_s2_byteenable),                   //       .byteenable
		.clk2        (parameter_clk_clk),                                //   clk2.clk
		.reset2      (rst_controller_001_reset_out_reset),               // reset2.reset
		.reset_req2  (rst_controller_001_reset_out_reset_req),           //       .reset_req
		.freeze      (1'b0)                                              // (terminated)
	);

	Pararameter_Comms_SYS_Reset reset (
		.clk        (pheriphal_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_reset_s1_readdata),   //                    .readdata
		.out_port   (reset_out_export)                       // external_connection.export
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (15),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge_0 (
		.m0_clk           (pheriphal_clk_clk),                           //   m0_clk.clk
		.m0_reset         (rst_controller_reset_out_reset),              // m0_reset.reset
		.s0_clk           (slave_clk_clk),                               //   s0_clk.clk
		.s0_reset         (slave_reset_reset),                           // s0_reset.reset
		.s0_waitrequest   (mapped_slave_waitrequest),                    //       s0.waitrequest
		.s0_readdata      (mapped_slave_readdata),                       //         .readdata
		.s0_readdatavalid (mapped_slave_readdatavalid),                  //         .readdatavalid
		.s0_burstcount    (mapped_slave_burstcount),                     //         .burstcount
		.s0_writedata     (mapped_slave_writedata),                      //         .writedata
		.s0_address       (mapped_slave_address),                        //         .address
		.s0_write         (mapped_slave_write),                          //         .write
		.s0_read          (mapped_slave_read),                           //         .read
		.s0_byteenable    (mapped_slave_byteenable),                     //         .byteenable
		.s0_debugaccess   (mapped_slave_debugaccess),                    //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_0_m0_waitrequest),   //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_0_m0_readdata),      //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_0_m0_readdatavalid), //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_0_m0_burstcount),    //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_0_m0_writedata),     //         .writedata
		.m0_address       (mm_clock_crossing_bridge_0_m0_address),       //         .address
		.m0_write         (mm_clock_crossing_bridge_0_m0_write),         //         .write
		.m0_read          (mm_clock_crossing_bridge_0_m0_read),          //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_0_m0_byteenable),    //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_0_m0_debugaccess)    //         .debugaccess
	);

	Pararameter_Comms_SYS_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                                   (pheriphal_clk_clk),                                //                                                 clk_0_clk.clk
		.mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                   // mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_0_m0_address                           (mm_clock_crossing_bridge_0_m0_address),            //                             mm_clock_crossing_bridge_0_m0.address
		.mm_clock_crossing_bridge_0_m0_waitrequest                       (mm_clock_crossing_bridge_0_m0_waitrequest),        //                                                          .waitrequest
		.mm_clock_crossing_bridge_0_m0_burstcount                        (mm_clock_crossing_bridge_0_m0_burstcount),         //                                                          .burstcount
		.mm_clock_crossing_bridge_0_m0_byteenable                        (mm_clock_crossing_bridge_0_m0_byteenable),         //                                                          .byteenable
		.mm_clock_crossing_bridge_0_m0_read                              (mm_clock_crossing_bridge_0_m0_read),               //                                                          .read
		.mm_clock_crossing_bridge_0_m0_readdata                          (mm_clock_crossing_bridge_0_m0_readdata),           //                                                          .readdata
		.mm_clock_crossing_bridge_0_m0_readdatavalid                     (mm_clock_crossing_bridge_0_m0_readdatavalid),      //                                                          .readdatavalid
		.mm_clock_crossing_bridge_0_m0_write                             (mm_clock_crossing_bridge_0_m0_write),              //                                                          .write
		.mm_clock_crossing_bridge_0_m0_writedata                         (mm_clock_crossing_bridge_0_m0_writedata),          //                                                          .writedata
		.mm_clock_crossing_bridge_0_m0_debugaccess                       (mm_clock_crossing_bridge_0_m0_debugaccess),        //                                                          .debugaccess
		.Parameter_GPIO_s1_address                                       (mm_interconnect_0_parameter_gpio_s1_address),      //                                         Parameter_GPIO_s1.address
		.Parameter_GPIO_s1_write                                         (mm_interconnect_0_parameter_gpio_s1_write),        //                                                          .write
		.Parameter_GPIO_s1_readdata                                      (mm_interconnect_0_parameter_gpio_s1_readdata),     //                                                          .readdata
		.Parameter_GPIO_s1_writedata                                     (mm_interconnect_0_parameter_gpio_s1_writedata),    //                                                          .writedata
		.Parameter_GPIO_s1_chipselect                                    (mm_interconnect_0_parameter_gpio_s1_chipselect),   //                                                          .chipselect
		.Parameter_RX_RAM_s1_address                                     (mm_interconnect_0_parameter_rx_ram_s1_address),    //                                       Parameter_RX_RAM_s1.address
		.Parameter_RX_RAM_s1_write                                       (mm_interconnect_0_parameter_rx_ram_s1_write),      //                                                          .write
		.Parameter_RX_RAM_s1_readdata                                    (mm_interconnect_0_parameter_rx_ram_s1_readdata),   //                                                          .readdata
		.Parameter_RX_RAM_s1_writedata                                   (mm_interconnect_0_parameter_rx_ram_s1_writedata),  //                                                          .writedata
		.Parameter_RX_RAM_s1_byteenable                                  (mm_interconnect_0_parameter_rx_ram_s1_byteenable), //                                                          .byteenable
		.Parameter_RX_RAM_s1_chipselect                                  (mm_interconnect_0_parameter_rx_ram_s1_chipselect), //                                                          .chipselect
		.Parameter_RX_RAM_s1_clken                                       (mm_interconnect_0_parameter_rx_ram_s1_clken),      //                                                          .clken
		.Parameter_TX_RAM_s1_address                                     (mm_interconnect_0_parameter_tx_ram_s1_address),    //                                       Parameter_TX_RAM_s1.address
		.Parameter_TX_RAM_s1_write                                       (mm_interconnect_0_parameter_tx_ram_s1_write),      //                                                          .write
		.Parameter_TX_RAM_s1_readdata                                    (mm_interconnect_0_parameter_tx_ram_s1_readdata),   //                                                          .readdata
		.Parameter_TX_RAM_s1_writedata                                   (mm_interconnect_0_parameter_tx_ram_s1_writedata),  //                                                          .writedata
		.Parameter_TX_RAM_s1_byteenable                                  (mm_interconnect_0_parameter_tx_ram_s1_byteenable), //                                                          .byteenable
		.Parameter_TX_RAM_s1_chipselect                                  (mm_interconnect_0_parameter_tx_ram_s1_chipselect), //                                                          .chipselect
		.Parameter_TX_RAM_s1_clken                                       (mm_interconnect_0_parameter_tx_ram_s1_clken),      //                                                          .clken
		.Reset_s1_address                                                (mm_interconnect_0_reset_s1_address),               //                                                  Reset_s1.address
		.Reset_s1_write                                                  (mm_interconnect_0_reset_s1_write),                 //                                                          .write
		.Reset_s1_readdata                                               (mm_interconnect_0_reset_s1_readdata),              //                                                          .readdata
		.Reset_s1_writedata                                              (mm_interconnect_0_reset_s1_writedata),             //                                                          .writedata
		.Reset_s1_chipselect                                             (mm_interconnect_0_reset_s1_chipselect)             //                                                          .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~pheriphal_reset_reset_n),           // reset_in0.reset
		.clk            (pheriphal_clk_clk),                  //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~parameter_reset_reset_n),               // reset_in0.reset
		.clk            (parameter_clk_clk),                      //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
