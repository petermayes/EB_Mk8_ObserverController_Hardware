// subsystemA.v

// Generated using ACDS version 18.1 646

`timescale 1 ps / 1 ps
module subsystemA (
		output wire [7:0]  led_gpio_external_connection_export, // led_gpio_external_connection.export
		output wire        mapped_slave_waitrequest,            //                 mapped_slave.waitrequest
		output wire [31:0] mapped_slave_readdata,               //                             .readdata
		output wire        mapped_slave_readdatavalid,          //                             .readdatavalid
		input  wire [0:0]  mapped_slave_burstcount,             //                             .burstcount
		input  wire [31:0] mapped_slave_writedata,              //                             .writedata
		input  wire [9:0]  mapped_slave_address,                //                             .address
		input  wire        mapped_slave_write,                  //                             .write
		input  wire        mapped_slave_read,                   //                             .read
		input  wire [3:0]  mapped_slave_byteenable,             //                             .byteenable
		input  wire        mapped_slave_debugaccess,            //                             .debugaccess
		input  wire        pheriphal_clk_clk,                   //                pheriphal_clk.clk
		input  wire        pheriphal_reset_reset_n,             //              pheriphal_reset.reset_n
		input  wire        slave_clk_clk,                       //                    slave_clk.clk
		input  wire        slave_reset_reset,                   //                  slave_reset.reset
		output wire [7:0]  tp_gpio_external_connection_export   //  tp_gpio_external_connection.export
	);

	wire         mm_clock_crossing_bridge_0_m0_waitrequest;   // mm_interconnect_0:mm_clock_crossing_bridge_0_m0_waitrequest -> mm_clock_crossing_bridge_0:m0_waitrequest
	wire  [31:0] mm_clock_crossing_bridge_0_m0_readdata;      // mm_interconnect_0:mm_clock_crossing_bridge_0_m0_readdata -> mm_clock_crossing_bridge_0:m0_readdata
	wire         mm_clock_crossing_bridge_0_m0_debugaccess;   // mm_clock_crossing_bridge_0:m0_debugaccess -> mm_interconnect_0:mm_clock_crossing_bridge_0_m0_debugaccess
	wire   [9:0] mm_clock_crossing_bridge_0_m0_address;       // mm_clock_crossing_bridge_0:m0_address -> mm_interconnect_0:mm_clock_crossing_bridge_0_m0_address
	wire         mm_clock_crossing_bridge_0_m0_read;          // mm_clock_crossing_bridge_0:m0_read -> mm_interconnect_0:mm_clock_crossing_bridge_0_m0_read
	wire   [3:0] mm_clock_crossing_bridge_0_m0_byteenable;    // mm_clock_crossing_bridge_0:m0_byteenable -> mm_interconnect_0:mm_clock_crossing_bridge_0_m0_byteenable
	wire         mm_clock_crossing_bridge_0_m0_readdatavalid; // mm_interconnect_0:mm_clock_crossing_bridge_0_m0_readdatavalid -> mm_clock_crossing_bridge_0:m0_readdatavalid
	wire  [31:0] mm_clock_crossing_bridge_0_m0_writedata;     // mm_clock_crossing_bridge_0:m0_writedata -> mm_interconnect_0:mm_clock_crossing_bridge_0_m0_writedata
	wire         mm_clock_crossing_bridge_0_m0_write;         // mm_clock_crossing_bridge_0:m0_write -> mm_interconnect_0:mm_clock_crossing_bridge_0_m0_write
	wire   [0:0] mm_clock_crossing_bridge_0_m0_burstcount;    // mm_clock_crossing_bridge_0:m0_burstcount -> mm_interconnect_0:mm_clock_crossing_bridge_0_m0_burstcount
	wire         mm_interconnect_0_tp_gpio_s1_chipselect;     // mm_interconnect_0:TP_GPIO_s1_chipselect -> TP_GPIO:chipselect
	wire  [31:0] mm_interconnect_0_tp_gpio_s1_readdata;       // TP_GPIO:readdata -> mm_interconnect_0:TP_GPIO_s1_readdata
	wire   [2:0] mm_interconnect_0_tp_gpio_s1_address;        // mm_interconnect_0:TP_GPIO_s1_address -> TP_GPIO:address
	wire         mm_interconnect_0_tp_gpio_s1_write;          // mm_interconnect_0:TP_GPIO_s1_write -> TP_GPIO:write_n
	wire  [31:0] mm_interconnect_0_tp_gpio_s1_writedata;      // mm_interconnect_0:TP_GPIO_s1_writedata -> TP_GPIO:writedata
	wire         mm_interconnect_0_led_gpio_s1_chipselect;    // mm_interconnect_0:LED_GPIO_s1_chipselect -> LED_GPIO:chipselect
	wire  [31:0] mm_interconnect_0_led_gpio_s1_readdata;      // LED_GPIO:readdata -> mm_interconnect_0:LED_GPIO_s1_readdata
	wire   [2:0] mm_interconnect_0_led_gpio_s1_address;       // mm_interconnect_0:LED_GPIO_s1_address -> LED_GPIO:address
	wire         mm_interconnect_0_led_gpio_s1_write;         // mm_interconnect_0:LED_GPIO_s1_write -> LED_GPIO:write_n
	wire  [31:0] mm_interconnect_0_led_gpio_s1_writedata;     // mm_interconnect_0:LED_GPIO_s1_writedata -> LED_GPIO:writedata
	wire         rst_controller_reset_out_reset;              // rst_controller:reset_out -> [LED_GPIO:reset_n, TP_GPIO:reset_n, mm_clock_crossing_bridge_0:m0_reset, mm_interconnect_0:mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset_reset]

	subsystemA_LED_GPIO led_gpio (
		.clk        (pheriphal_clk_clk),                        //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_led_gpio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_gpio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_gpio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_gpio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_gpio_s1_readdata),   //                    .readdata
		.out_port   (led_gpio_external_connection_export)       // external_connection.export
	);

	subsystemA_LED_GPIO tp_gpio (
		.clk        (pheriphal_clk_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_tp_gpio_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_tp_gpio_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_tp_gpio_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_tp_gpio_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_tp_gpio_s1_readdata),   //                    .readdata
		.out_port   (tp_gpio_external_connection_export)       // external_connection.export
	);

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.HDL_ADDR_WIDTH      (10),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (4),
		.RESPONSE_FIFO_DEPTH (4),
		.MASTER_SYNC_DEPTH   (2),
		.SLAVE_SYNC_DEPTH    (2)
	) mm_clock_crossing_bridge_0 (
		.m0_clk           (pheriphal_clk_clk),                           //   m0_clk.clk
		.m0_reset         (rst_controller_reset_out_reset),              // m0_reset.reset
		.s0_clk           (slave_clk_clk),                               //   s0_clk.clk
		.s0_reset         (slave_reset_reset),                           // s0_reset.reset
		.s0_waitrequest   (mapped_slave_waitrequest),                    //       s0.waitrequest
		.s0_readdata      (mapped_slave_readdata),                       //         .readdata
		.s0_readdatavalid (mapped_slave_readdatavalid),                  //         .readdatavalid
		.s0_burstcount    (mapped_slave_burstcount),                     //         .burstcount
		.s0_writedata     (mapped_slave_writedata),                      //         .writedata
		.s0_address       (mapped_slave_address),                        //         .address
		.s0_write         (mapped_slave_write),                          //         .write
		.s0_read          (mapped_slave_read),                           //         .read
		.s0_byteenable    (mapped_slave_byteenable),                     //         .byteenable
		.s0_debugaccess   (mapped_slave_debugaccess),                    //         .debugaccess
		.m0_waitrequest   (mm_clock_crossing_bridge_0_m0_waitrequest),   //       m0.waitrequest
		.m0_readdata      (mm_clock_crossing_bridge_0_m0_readdata),      //         .readdata
		.m0_readdatavalid (mm_clock_crossing_bridge_0_m0_readdatavalid), //         .readdatavalid
		.m0_burstcount    (mm_clock_crossing_bridge_0_m0_burstcount),    //         .burstcount
		.m0_writedata     (mm_clock_crossing_bridge_0_m0_writedata),     //         .writedata
		.m0_address       (mm_clock_crossing_bridge_0_m0_address),       //         .address
		.m0_write         (mm_clock_crossing_bridge_0_m0_write),         //         .write
		.m0_read          (mm_clock_crossing_bridge_0_m0_read),          //         .read
		.m0_byteenable    (mm_clock_crossing_bridge_0_m0_byteenable),    //         .byteenable
		.m0_debugaccess   (mm_clock_crossing_bridge_0_m0_debugaccess)    //         .debugaccess
	);

	subsystemA_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                                   (pheriphal_clk_clk),                           //                                                 clk_0_clk.clk
		.mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),              // mm_clock_crossing_bridge_0_m0_reset_reset_bridge_in_reset.reset
		.mm_clock_crossing_bridge_0_m0_address                           (mm_clock_crossing_bridge_0_m0_address),       //                             mm_clock_crossing_bridge_0_m0.address
		.mm_clock_crossing_bridge_0_m0_waitrequest                       (mm_clock_crossing_bridge_0_m0_waitrequest),   //                                                          .waitrequest
		.mm_clock_crossing_bridge_0_m0_burstcount                        (mm_clock_crossing_bridge_0_m0_burstcount),    //                                                          .burstcount
		.mm_clock_crossing_bridge_0_m0_byteenable                        (mm_clock_crossing_bridge_0_m0_byteenable),    //                                                          .byteenable
		.mm_clock_crossing_bridge_0_m0_read                              (mm_clock_crossing_bridge_0_m0_read),          //                                                          .read
		.mm_clock_crossing_bridge_0_m0_readdata                          (mm_clock_crossing_bridge_0_m0_readdata),      //                                                          .readdata
		.mm_clock_crossing_bridge_0_m0_readdatavalid                     (mm_clock_crossing_bridge_0_m0_readdatavalid), //                                                          .readdatavalid
		.mm_clock_crossing_bridge_0_m0_write                             (mm_clock_crossing_bridge_0_m0_write),         //                                                          .write
		.mm_clock_crossing_bridge_0_m0_writedata                         (mm_clock_crossing_bridge_0_m0_writedata),     //                                                          .writedata
		.mm_clock_crossing_bridge_0_m0_debugaccess                       (mm_clock_crossing_bridge_0_m0_debugaccess),   //                                                          .debugaccess
		.LED_GPIO_s1_address                                             (mm_interconnect_0_led_gpio_s1_address),       //                                               LED_GPIO_s1.address
		.LED_GPIO_s1_write                                               (mm_interconnect_0_led_gpio_s1_write),         //                                                          .write
		.LED_GPIO_s1_readdata                                            (mm_interconnect_0_led_gpio_s1_readdata),      //                                                          .readdata
		.LED_GPIO_s1_writedata                                           (mm_interconnect_0_led_gpio_s1_writedata),     //                                                          .writedata
		.LED_GPIO_s1_chipselect                                          (mm_interconnect_0_led_gpio_s1_chipselect),    //                                                          .chipselect
		.TP_GPIO_s1_address                                              (mm_interconnect_0_tp_gpio_s1_address),        //                                                TP_GPIO_s1.address
		.TP_GPIO_s1_write                                                (mm_interconnect_0_tp_gpio_s1_write),          //                                                          .write
		.TP_GPIO_s1_readdata                                             (mm_interconnect_0_tp_gpio_s1_readdata),       //                                                          .readdata
		.TP_GPIO_s1_writedata                                            (mm_interconnect_0_tp_gpio_s1_writedata),      //                                                          .writedata
		.TP_GPIO_s1_chipselect                                           (mm_interconnect_0_tp_gpio_s1_chipselect)      //                                                          .chipselect
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~pheriphal_reset_reset_n),       // reset_in0.reset
		.clk            (pheriphal_clk_clk),              //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
